//////////////////////////////////////////////////////////////////////////////////
// Test bench for Exercise #9  
// Student Name:
// Date: 
//
// Description: A testbench module to test Ex9
// You need to write the whole file
//////////////////////////////////////////////////////////////////////////////////

